library IEEE;
use IEEE.std_logic_1164.all  ; 
use IEEE.std_logic_arith.all  ; 
use IEEE.std_logic_unsigned.all  ; 
entity testbench is
end entity;

architecture arc of testbench is
	constant not_data_constant:std_logic_vector:="000000000000000000000011010111101111100110110110011011111001101111110011011110001101101100110111100011011011110101111100110101111110101010011110000000000000000000000000000000000000000011010111110111110011011011001101111100110111110011011110001101101100011011110001101101111010111110011010111110101010011110000000000000000000000000000000000000000000000000000000001101011110111110011011011001100111110011011111001101111000110110110011011110001101101111011011111001101011111010101001111000000000000000000000000000000000000000001101011110111110011011011001101111100110111110011011110000110110110011011110001101101111010111110011010111110101010001111000000000000000000000000000000000011010111101111100110110110011011111001101111100110111100001101101100110111100011011011110101111100110101111101010100011110000000000000000000000000000000000000110101111011111001101100110011011111001101111100110111100011011011001101111000110111011110101111100110101111101010100111100000000000000000000000000000110101111011111100110110110011011111001101111100110111100011011011001100111100011011011110101111100110101111101010100111100000000000000000000000000000000000000000000001101011110111110011011011001101111100111011111001101111000110110110011011110001101101111010111110001101011111010101001111000000000000000000000000000000000000000000000000000000000001101011110111110011011011001101111100110111111001101111000110110110011011110001101101111010111110011101011111010101001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101111011111100110110110011011111001101111100110111100011011011001100111100011011011110101111100110101111101010100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101111011111001101101100110111110001101111100110111100011011011001101111000110110111101011111100110101111101010100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100101111011111001101101100110111110011011111001101111000110111011001101111000110110111101011111001101011111010101001111000000000000000000000000000000000000000000011010111101111100110110110011101111100110111110011011110001101101100110111100011011011111010111110011010111110101010011110000000000000000";
	signal not_data:std_logic;
	signal successful:std_logic;
	signal ID:std_logic_vector(39 downto 0); 
	signal data:std_logic;
	signal reset:std_logic:='1';
		-- According to the communication protocol, the data
		-- being send are ASCII codes represnting the characters:
		-- [0-9] and [A-F]. There for the ASCII codes are:
		--   code[bin]   | code[dec] | character
		-- =====================================
		--   0b00011110  |    30     |    0
		--   0b00011111  |    31     |    1
		--   0b00100000  |    32     |    2
		--   0b00100001  |    33     |    3
		--   0b00100010  |    34     |    4
		--   0b00100011  |    35     |    5
		--   0b00100100  |    36     |    6
		--   0b00100101  |    37     |    7
		--   0b00100110  |    38     |    8
		--   0b00100111  |    39     |    9
		--   0b00101001  |    41     |    A
		--   0b00101010  |    42     |    B
		--   0b00101011  |    43     |    C
		--   0b00101100  |    44     |    D
		--   0b00101101  |    45     |    E
		--   0b00101110  |    46     |    F
		-- Therefor, the maximum number of zeros appears with 32[dec]
		-- - The longest sequence of zeros is of 5.
		-- If our sampling rate (for example) 16 times higher then
		-- Nyquist's minimum, then for a sequence of 5 zeros in the
		-- data stream we should count 5*16 samples of the same state.
		-- If 5*16=80 then we need ciel(log2(80))=7 bits for `samples`
		-- that's the minimal number of bits to represent the number 80.
	constant extra_samples_width:integer:=7;
	signal samples:std_logic_vector(extra_samples_width-1 downto 0);
	signal clk50mhz:std_logic:='0';
	signal PLL_clk:std_logic:='0';
	signal data_clk:std_logic:='0';
	component data_buffer
		generic(
			extra_samples_width:integer:=4
		);
		port(
			clk		:in std_logic;
			reset	:in std_logic;
			not_data:in std_logic;
			data	:out std_logic;
			samples	:out std_logic_vector(extra_samples_width-1 downto 0)
		);
	end component;
begin
	clk50mhz<=not clk50mhz after 10 ns;--10[ns]=(1/100mhz)/2,t(50mhz)=20ns
	reset<='0','1' after 1 us;
	PLL_clk<=not PLL_clk after 10 us;
	data_clk<=not data_clk after 160 us;
	data_buffer_inst:data_buffer
		generic map(
			extra_samples_width=>extra_samples_width
		)
		port map(
			clk		=>PLL_clk,
			reset	=>reset,
			not_data=>not_data,
			data	=>data,
			samples	=>samples
		);
	process(data_clk,reset)
		variable counter:integer;
	begin
		if reset='0' then
			counter:=0;
			not_data<='1';
		elsif rising_edge(data_clk) then
			counter:=counter+1;
			if counter<not_data_constant'length then
				not_data<=not_data_constant(counter);
			else
				counter:=0;
			end if;
		end if;
	end process;
end;
