library IEEE;
use IEEE.std_logic_1164.all  ; 
use IEEE.std_logic_arith.all  ; 
use IEEE.std_logic_unsigned.all  ; 
entity testbench is
end entity;

architecture arc of testbench is
	constant not_data_constant:std_logic_vector:="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110110011011111001101111110011011110001101101100110111100011011011110101111100110101111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111110111110011011011001101111100110111110011011110001101101100011011110001101101111010111110011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101011110111110011011011001100111110011011111001101111000110110110011011110001101101111011011111001101011111010101001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110110011011111001101111100110111100001101101100110111100011011011110101111100110101111101010100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110110011011111001101111100110111100001101101100110111100011011011110101111100110101111101010100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110011001101111100110111110011011110001101101100110111100011011101111010111110011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111110011011011001101111100110111110011011110001101101100110011110001101101111010111110011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110110011011111001110111110011011110001101101100110111100011011011110101111100011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101111011111001101101100110111110011011111100110111100011011011001101111000110110111101011111001110101111101010100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111110011011011001101111100110111110011011110001101101100110011110001101101111010111110011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110110011011111000110111110011011110001101101100110111100011011011110101111110011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010111101111100110110110011011111001101111100110111100011011101100110111100011011011110101111100110101111101010100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110110011101111100110111110011011110001101101100110111100011011011111010111110011010111110101010011110000000000000000";
	signal not_data:std_logic;
	signal successful:std_logic;
	signal ID:std_logic_vector(39 downto 0); 
	signal data:std_logic;
	signal reset:std_logic:='1';
	signal samples:std_logic_vector(15 downto 0);
	signal clk50mhz:std_logic:='0';
	signal PLL_clk:std_logic:='0';--clk2400hz 
	component data_buffer
		port(
			clk384000hz	:in std_logic;
			reset		:in std_logic;
			not_data	:in std_logic;
			data		:out std_logic;
			samples		:out std_logic_vector(15 downto 0)
		);
	end component;
begin
	clk50mhz<=not clk50mhz after 10 ns;--10[ns]=(1/100mhz)/2,t(50mhz)=20ns
	reset<='0','1' after 1 us;
	PLL_clk<=not PLL_clk after 2604 ns;--2604[ns]=(1/384000hz)
	data_buffer_inst:data_buffer
		port map(
			clk384000hz	=>PLL_clk,
			reset		=>reset,
			not_data	=>not_data,
			data		=>data,
			samples		=>samples
		);
	process(PLL_clk,reset)
		variable counter:integer;
	begin
		if reset='0' then
			counter:=0;
			not_data<='1';
		elsif rising_edge(PLL_clk) then
			counter:=counter+1;
			if (counter<not_data_constant'length)then
				not_data<=not_data_constant(not_data_constant'length-1);
			else
				counter:=0;
			end if;
		end if;
	end process;
end;
