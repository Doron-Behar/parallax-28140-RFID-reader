library IEEE;
use IEEE.std_logic_1164.all  ; 
use IEEE.std_logic_arith.all  ; 
use IEEE.std_logic_unsigned.all  ; 
entity testbench is
end entity;

architecture arc of testbench is
	constant not_data_constant:std_logic_vector:="00001101011110111110011011011001101111100110111111001101111000110110110011011110001101101111010111110011010111111010101001111000000000000110101111101111100110110110011011111001101111100110111100011011011000110111100011011011110101111100110101111101010100111100000000011010111101111100110110110011001111100110111110011011110001101101100110111100011011011110110111110011010111110101010011110000000000011010111101111100110110110011011111001101111100110111100001101101100110111100011011011110101111100110101111101010100011110000000000000110101111011111001101101100110111110011011111001101111000011011011001101111000110110111101011111001101011111010101000111100000000011010111101111100110110011001101111100110111110011011110001101101100110111100011011101111010111110011010111110101010011110000000000000011010111101111110011011011001101111100110111110011011110001101101100110011110001101101111010111110011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110110011011111001110111110011011110001101101100110111100011011011110101111100011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101111011111001101101100110111110011011111100110111100011011011001101111000110110111101011111001110101111101010100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111110011011011001101111100110111110011011110001101101100110011110001101101111010111110011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110110011011111000110111110011011110001101101100110111100011011011110101111110011010111110101010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010111101111100110110110011011111001101111100110111100011011101100110111100011011011110101111100110101111101010100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010111101111100110110110011101111100110111110011011110001101101100110111100011011011111010111110011010111110101010011110000000000000000";
	signal not_data:std_logic;
	signal successful:std_logic;
	signal ID:std_logic_vector(39 downto 0); 
	signal data:std_logic;
	signal reset:std_logic:='1';
	constant extra_samples_width:integer:=4;
	signal samples:std_logic_vector(extra_samples_width-1 downto 0);
	signal clk50mhz:std_logic:='0';
	signal PLL_clk:std_logic:='0';
	signal data_clk:std_logic:='0';
	component data_buffer
		generic(
			extra_samples_width:integer:=4
		);
		port(
			clk		:in std_logic;
			reset	:in std_logic;
			not_data:in std_logic;
			data	:out std_logic;
			samples	:out std_logic_vector(extra_samples_width-1 downto 0)
		);
	end component;
begin
	clk50mhz<=not clk50mhz after 10 ns;--10[ns]=(1/100mhz)/2,t(50mhz)=20ns
	reset<='0','1' after 1 us;
	PLL_clk<=not PLL_clk after 10 us;
	data_clk<=not data_clk after 80 us;
	data_buffer_inst:data_buffer
		generic map(
			extra_samples_width=>4
		)
		port map(
			clk		=>PLL_clk,
			reset	=>reset,
			not_data=>not_data,
			data	=>data,
			samples	=>samples
		);
	process(data_clk,reset)
		variable counter:integer;
	begin
		if reset='0' then
			counter:=0;
			not_data<='1';
		elsif rising_edge(data_clk) then
			counter:=counter+1;
			if counter<not_data_constant'length then
				not_data<=not_data_constant(counter);
			else
				counter:=0;
			end if;
		end if;
	end process;
end;
